`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/11/30 15:19:44
// Design Name: 
// Module Name: backgroundcolor_map
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module backgroundcolor_map(  input logic[7:0] background_red,
                                output logic[23:0] background_rgb
        

    );
    always_comb begin
        unique case(background_red)
            8'h88: background_rgb=24'h889166;
            8'h82: background_rgb=24'h828b5e;
            8'h95: background_rgb=24'h95a16b;
            8'h48: background_rgb=24'h484939;
            8'h00: background_rgb=24'h000000;
            8'h84: background_rgb=24'h848d5f;
            8'h91: background_rgb=24'h919c68;
            8'h34: background_rgb=24'h34322c;
            8'h46: background_rgb=24'h464638;
            8'h8f: background_rgb=24'h8f9a67;
            8'h70: background_rgb=24'h707652;
            8'h1c: background_rgb=24'h1c161d;
            8'h85: background_rgb=24'h858f60;
            8'h87: background_rgb=24'h879162;
            8'h56: background_rgb=24'h565942;
            8'h3a: background_rgb=24'h3a3830;
            8'h93: background_rgb=24'h939e6a;
            8'h83: background_rgb=24'h838c5f;
            8'h8d: background_rgb=24'h8d9766;
            8'h2e: background_rgb=24'h2e2b29;
            8'h2f: background_rgb=24'h2f2d26;
            8'h6f: background_rgb=24'h6f7a49;
            8'h64: background_rgb=24'h646c42;
            8'h62: background_rgb=24'h626b42;
            8'h71: background_rgb=24'h717c4a;
            8'h3b: background_rgb=24'h3b3b2c;
            8'h37: background_rgb=24'h37372a;
            8'h6d: background_rgb=24'h6d7647;
            8'h55: background_rgb=24'h555b3b;
            8'h03: background_rgb=24'h03000d;
            8'h19: background_rgb=24'h19131a;
            8'h65: background_rgb=24'h656d43;
            8'h66: background_rgb=24'h667044;
            8'h6b: background_rgb=24'h6b7446;
            8'h23: background_rgb=24'h231f1f;
            8'h4e: background_rgb=24'h4e3432;
            8'h76: background_rgb=24'h765044;
            8'h4f: background_rgb=24'h4f3432;
            8'h49: background_rgb=24'h49312a;
            8'hbf: background_rgb=24'hbf8655;
            8'ha9: background_rgb=24'ha9774e;
            8'hba: background_rgb=24'hba8354;
            8'h90: background_rgb=24'h906544;
            8'h1a: background_rgb=24'h1a171d;
            8'h39: background_rgb=24'h39323a;
            8'h98: background_rgb=24'h989390;
            8'h79: background_rgb=24'h797374;
            8'h0d: background_rgb=24'h0d0315;
            8'h16: background_rgb=24'h160d17;
            8'h60: background_rgb=24'h607490;
            8'ha7: background_rgb=24'ha7d6ff;
            8'h9b: background_rgb=24'h9bc6ed;
            8'h89: background_rgb=24'h89acd1;
            8'h0e: background_rgb=24'h0e071b;
            8'h0c: background_rgb=24'h0c0108;
            8'h7b: background_rgb=24'h7b835a;
            8'h8b: background_rgb=24'h8b9665;
            8'h43: background_rgb=24'h434531;
            8'h09: background_rgb=24'h090011;
            8'h21: background_rgb=24'h211b20;
            8'h1e: background_rgb=24'h1e181e;
            8'h69: background_rgb=24'h697346;
            8'h5d: background_rgb=24'h5d653f;
            8'h0b: background_rgb=24'h0b0211;
            8'h10: background_rgb=24'h100716;
            8'h4b: background_rgb=24'h4b4c3b;
            8'h96: background_rgb=24'h96a26c;
            8'h8a: background_rgb=24'h8a9564;
            8'h7d: background_rgb=24'h7d855b;
            8'h12: background_rgb=24'h120917;
            8'h5c: background_rgb=24'h5c643f;
            8'h6a: background_rgb=24'h6a7346;
            8'h63: background_rgb=24'h636b42;
            8'h57: background_rgb=24'h575e3c;
            8'h25: background_rgb=24'h252822;
            8'h27: background_rgb=24'h272a23;
            8'h29: background_rgb=24'h292c24;
            8'h2b: background_rgb=24'h2b2f25;
            8'h5f: background_rgb=24'h5f6640;
            8'h68: background_rgb=24'h687145;
            8'h44: background_rgb=24'h44453f;
            8'h47: background_rgb=24'h474841;
            8'h2d: background_rgb=24'h2d2c30;
            8'h38: background_rgb=24'h383738;
            8'h41: background_rgb=24'h41423e;
            8'h30: background_rgb=24'h302d33;
            8'h35: background_rgb=24'h353336;
            8'h45: background_rgb=24'h454540;
            8'h3d: background_rgb=24'h3d3d3b;
            8'h3f: background_rgb=24'h3f403b;
            8'h31: background_rgb=24'h312e33;
            8'h40: background_rgb=24'h40403b;
            8'h36: background_rgb=24'h363436;
            8'h3c: background_rgb=24'h3c3739;
            8'h42: background_rgb=24'h423c3c;
            8'h4d: background_rgb=24'h4d443e;
            8'h4a: background_rgb=24'h4a413d;
            8'h4c: background_rgb=24'h4c433e;
            8'h32: background_rgb=24'h323034;
            8'h33: background_rgb=24'h333135;
            8'h3e: background_rgb=24'h3e3f3b;
            8'h28: background_rgb=24'h282b24;
            8'h2a: background_rgb=24'h2a2c22;
            8'h2c: background_rgb=24'h2c2932;
            8'h1f: background_rgb=24'h1f231c;
            8'h22: background_rgb=24'h222420;
            8'h24: background_rgb=24'h242721;
            8'h26: background_rgb=24'h262a20;
            8'ha3: background_rgb=24'ha3a099;
            8'h9e: background_rgb=24'h9e9b94;
            8'ha1: background_rgb=24'ha19f98;
            8'hb6: background_rgb=24'hb6b3ab;
            8'hb7: background_rgb=24'hb7b3ac;
            8'hb8: background_rgb=24'hb8b4ad;
            8'ha4: background_rgb=24'ha4a19a;
            8'h9a: background_rgb=24'h9a9891;
            8'ha6: background_rgb=24'ha6a39c;
            8'h7a: background_rgb=24'h7a7677;
            8'haa: background_rgb=24'haaa8a8;
            8'h6c: background_rgb=24'h6c6768;
            8'h9c: background_rgb=24'h9c9992;
            8'hbe: background_rgb=24'hbebbb4;
            8'hb2: background_rgb=24'hb2aea7;
            8'h1d: background_rgb=24'h1d201b;
            8'h73: background_rgb=24'h73726c;
            8'hb1: background_rgb=24'hb1aea6;
            8'hd4: background_rgb=24'hd4d0c6;
            8'hd2: background_rgb=24'hd2cec3;
            8'hd9: background_rgb=24'hd9d6ca;
            8'hc7: background_rgb=24'hc7c4b9;
            8'h8e: background_rgb=24'h8e8d82;
            8'h8c: background_rgb=24'h8c8c81;
            8'hc0: background_rgb=24'hc0bdb2;
            8'hdb: background_rgb=24'hdbd8cc;
            8'hcf: background_rgb=24'hcfccc0;
            8'hd7: background_rgb=24'hd7d4c7;
            8'hf0: background_rgb=24'hf0edde;
            8'hd5: background_rgb=24'hd5d2c6;
            8'h7c: background_rgb=24'h7c7575;
            8'he4: background_rgb=24'he4e2e1;
            8'hbd: background_rgb=24'hbdb9b8;
            8'h80: background_rgb=24'h807979;
            8'hd6: background_rgb=24'hd6d3c7;
            8'h86: background_rgb=24'h86867b;
            8'h20: background_rgb=24'h20241c;
            8'hef: background_rgb=24'hefebde;
            8'hc2: background_rgb=24'hc2bfb6;
            8'hc1: background_rgb=24'hc1beb4;
            8'hd8: background_rgb=24'hd8d5cb;
            8'h13: background_rgb=24'h13170f;
            8'h02: background_rgb=24'h020600;
            8'h94: background_rgb=24'h949289;
            8'hde: background_rgb=24'hded9cf;
            8'h7e: background_rgb=24'h7e7878;
            8'h74: background_rgb=24'h746e6e;
            8'had: background_rgb=24'hada9a9;
            8'h77: background_rgb=24'h777171;
            8'hcc: background_rgb=24'hccc9bf;
            8'h05: background_rgb=24'h050a02;
            8'hc5: background_rgb=24'hc5c1b7;
            8'hdf: background_rgb=24'hdfdcd1;
            8'ha0: background_rgb=24'ha09d94;
            8'hca: background_rgb=24'hcac7bd;
            8'hb9: background_rgb=24'hb9b6ac;
            8'h1b: background_rgb=24'h1b1f17;
            8'hbb: background_rgb=24'hbbb8af;
            8'hf6: background_rgb=24'hf6f3e4;
            8'h06: background_rgb=24'h06060b;
            8'h7f: background_rgb=24'h7f7a7a;
            8'hdd: background_rgb=24'hdddcdc;
            8'hb5: background_rgb=24'hb5b1b1;
            8'h18: background_rgb=24'h181c14;
            8'h92: background_rgb=24'h929087;
            8'hc9: background_rgb=24'hc9c6bb;
            8'h59: background_rgb=24'h595657;
            8'h81: background_rgb=24'h817b7b;
            8'h9d: background_rgb=24'h9d9999;
            8'h0f: background_rgb=24'h0f130c;
            8'h97: background_rgb=24'h97958c;
            8'hda: background_rgb=24'hdad7ca;
            8'hac: background_rgb=24'haca7a7;
            8'he1: background_rgb=24'he1e0e0;
            8'hb0: background_rgb=24'hb0acac;
            8'hbc: background_rgb=24'hbcb9b0;
            8'hc3: background_rgb=24'hc3c0b6;
            8'hd3: background_rgb=24'hd3cfc5;
            8'hdc: background_rgb=24'hdcd9cc;
            8'hf1: background_rgb=24'hf1eedf;
            8'h15: background_rgb=24'h15151a;
            8'h51: background_rgb=24'h514e51;
            8'h75: background_rgb=24'h756e6e;
            8'h58: background_rgb=24'h585951;
            8'hae: background_rgb=24'haeaba3;
            8'h52: background_rgb=24'h524f51;
            8'h04: background_rgb=24'h040801;
            8'h08: background_rgb=24'h080c04;
            8'h11: background_rgb=24'h111016;
            8'h53: background_rgb=24'h535051;
            8'hf7: background_rgb=24'hf7f4e6;
            8'hcb: background_rgb=24'hcbc8bd;
            8'hec: background_rgb=24'hece9db;
            8'hb3: background_rgb=24'hb3b0a7;
            8'hc4: background_rgb=24'hc4c1b7;
            8'h67: background_rgb=24'h676363;
            8'he3: background_rgb=24'he3e1d2;
            8'h72: background_rgb=24'h726c6d;
            8'hff: background_rgb=24'hffff58;
            8'hc6: background_rgb=24'hc6c3b7;
            8'hce: background_rgb=24'hcecbbf;
            8'h0a: background_rgb=24'h0a0a0f;
            8'hd0: background_rgb=24'hd0cdc1;
            8'he2: background_rgb=24'he2dfd2;
            8'h6e: background_rgb=24'h6e6e65;
            8'hcd: background_rgb=24'hcdcabe;
            8'h5a: background_rgb=24'h5a5856;
            8'he8: background_rgb=24'he8e7d6;
            8'hf4: background_rgb=24'hf4ce49;
            8'haf: background_rgb=24'hafaca3;
            8'he0: background_rgb=24'he0dcd2;
            8'h61: background_rgb=24'h615026;
            8'hd1: background_rgb=24'hd1cec1;
            8'h5e: background_rgb=24'h5e5c5b;
            8'hab: background_rgb=24'haba9a0;
            8'hc8: background_rgb=24'hc8a73f;
            8'hfa: background_rgb=24'hfaf8e6;
            8'h99: background_rgb=24'h99832d;
            8'hb4: background_rgb=24'hb48841;
            8'ha8: background_rgb=24'ha8a59e;
            8'ha5: background_rgb=24'ha58b36;
            8'hf2: background_rgb=24'hf2d349;
            8'he9: background_rgb=24'he9e5da;
            8'h5b: background_rgb=24'h5b5a59;
            8'he5: background_rgb=24'he5e0d5;
            8'hf3: background_rgb=24'hf3f1df;
            8'hee: background_rgb=24'heecc45;
            8'hf8: background_rgb=24'hf8d849;
            8'h54: background_rgb=24'h544e52;
            8'hed: background_rgb=24'hedecda;
            8'he7: background_rgb=24'he7cc48;
            8'h9f: background_rgb=24'h9f9b9b;
            8'h78: background_rgb=24'h787171;
            8'hfd: background_rgb=24'hfddc47;
            8'he6: background_rgb=24'he6b54b;
            8'hfe: background_rgb=24'hfec853;
            8'heb: background_rgb=24'hebe6da;
            8'hfb: background_rgb=24'hfbc650;
            8'h14: background_rgb=24'h140b16;
            8'hf5: background_rgb=24'hf5f1e4;
            8'h50: background_rgb=24'h505249;
            8'hf9: background_rgb=24'hf9f3e8;
            8'h07: background_rgb=24'h070b05;
            8'hea: background_rgb=24'heab94d;
            8'h17: background_rgb=24'h171a12;
            8'ha2: background_rgb=24'ha27e3a;
            8'h01: background_rgb=24'h010500;

        endcase
    end
endmodule
