`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/11/05 23:00:06
// Design Name: 
// Module Name: joeinstance
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
// the module is used to check whether the point is in square of center

module joe_color(  input logic[7:0] joe_red,
                   output logic[23:0] joe_rgb

    );
    always_comb 
    begin
    unique case(joe_red)
    8'hff: joe_rgb=24'hffffff;
    8'hc3: joe_rgb=24'hc37a78;
    8'h95: joe_rgb=24'h951211;
    8'ha4: joe_rgb=24'ha42928;
    8'ha3: joe_rgb=24'ha32422;
    8'h97: joe_rgb=24'h971615;
    8'hde: joe_rgb=24'hdec3c2;
    8'hc1: joe_rgb=24'hc17773;
    8'h8b: joe_rgb=24'h8b0000;
    8'h9d: joe_rgb=24'h9d110f;
    8'h9c: joe_rgb=24'h9c0908;
    8'h8e: joe_rgb=24'h8e0000;
    8'he0: joe_rgb=24'he0d4d0;
    8'hf3: joe_rgb=24'hf3ebea;
    8'hb7: joe_rgb=24'hb76f6b;
    8'hb9: joe_rgb=24'hb96f6b;
    8'ha8: joe_rgb=24'ha83936;
    8'h99: joe_rgb=24'h990a09;
    8'h9e: joe_rgb=24'h9e1513;
    8'h9b: joe_rgb=24'h9b0e0c;
    8'hb1: joe_rgb=24'hb15a56;
    8'hb2: joe_rgb=24'hb26460;
    8'hcb: joe_rgb=24'hcb9d99;
    8'hef: joe_rgb=24'hefe0df;
    8'ha0: joe_rgb=24'ha01916;
    8'h9f: joe_rgb=24'h9f1512;
    8'h82: joe_rgb=24'h820000;
    8'ha7: joe_rgb=24'ha7423f;
    8'hf7: joe_rgb=24'hf7f8f7;
    8'h9a: joe_rgb=24'h9a1412;
    8'h92: joe_rgb=24'h920000;
    8'hb4: joe_rgb=24'hb46360;
    8'hfe: joe_rgb=24'hfefdfc;
    8'hfd: joe_rgb=24'hfdfcfa;
    8'hfc: joe_rgb=24'hfcfaf8;
    8'hfa: joe_rgb=24'hfaf8f4;
    8'hfb: joe_rgb=24'hfbf9f5;
    8'hf5: joe_rgb=24'hf5f4f2;
    8'hb6: joe_rgb=24'hb66764;
    8'hb3: joe_rgb=24'hb35451;
    8'hb0: joe_rgb=24'hb04140;
    8'he6: joe_rgb=24'he6d978;
    8'hab: joe_rgb=24'hab3534;
    8'h93: joe_rgb=24'h930000;
    8'haa: joe_rgb=24'haa4b49;
    8'hd4: joe_rgb=24'hd4a7a4;
    8'ha1: joe_rgb=24'ha1700b;
    8'h96: joe_rgb=24'h965f05;
    8'hf0: joe_rgb=24'hf0efed;
    8'h90: joe_rgb=24'h900502;
    8'h8a: joe_rgb=24'h8a0000;
    8'h91: joe_rgb=24'h910000;
    8'h7e: joe_rgb=24'h7e0000;
    8'hb8: joe_rgb=24'hb85554;
    8'h7d: joe_rgb=24'h7d0000;
    8'hbe: joe_rgb=24'hbe6e6c;
    8'hac: joe_rgb=24'hac822a;
    8'hf2: joe_rgb=24'hf2f1ef;
    8'ha2: joe_rgb=24'ha21e1c;
    8'hb5: joe_rgb=24'hb54c4b;
    8'had: joe_rgb=24'had3b39;
    8'h8d: joe_rgb=24'h8d0000;
    8'hc6: joe_rgb=24'hc6817f;
    8'hee: joe_rgb=24'heee8da;
    8'hf9: joe_rgb=24'hf9f8f5;
    8'h8f: joe_rgb=24'h8f0000;
    8'hae: joe_rgb=24'hae3b3a;
    8'hc2: joe_rgb=24'hc29842;
    8'hba: joe_rgb=24'hba9242;
    8'ha9: joe_rgb=24'ha92f2e;
    8'hc7: joe_rgb=24'hc79d48;
    8'ha5: joe_rgb=24'ha57514;
    8'hf8: joe_rgb=24'hf8f6f3;
    8'hc4: joe_rgb=24'hc49a45;
    8'hf1: joe_rgb=24'hf1f0ee;
    8'h8c: joe_rgb=24'h8c0000;
    8'h94: joe_rgb=24'h940000;
    8'hc5: joe_rgb=24'hc57d7b;
    8'hc8: joe_rgb=24'hc89e49;
    8'h80: joe_rgb=24'h800000;
    8'hbf: joe_rgb=24'hbf7976;
    8'he2: joe_rgb=24'he2d0cd;
    8'hdf: joe_rgb=24'hdfcac7;
    8'hd6: joe_rgb=24'hd6b5b2;
    8'hdb: joe_rgb=24'hdbc1be;
    8'hed: joe_rgb=24'hede2e0;
    8'h81: joe_rgb=24'h810000;
    8'haf: joe_rgb=24'haf5450;
    8'hc9: joe_rgb=24'hc99794;
    8'h89: joe_rgb=24'h890000;
    8'h87: joe_rgb=24'h870000;
    8'h88: joe_rgb=24'h880000;
    8'he5: joe_rgb=24'he5d5d1;
    8'hd1: joe_rgb=24'hd1c3c0;
    8'h7a: joe_rgb=24'h7a6867;
    8'h71: joe_rgb=24'h715f60;
    8'he8: joe_rgb=24'he8dbd8;
    8'h66: joe_rgb=24'h666f6f;
    8'h5b: joe_rgb=24'h5b6467;
    8'ha6: joe_rgb=24'ha6781b;
    8'hda: joe_rgb=24'hdad3d0;
    8'hd5: joe_rgb=24'hd5b9a5;
    8'hec: joe_rgb=24'hecdac7;
    8'h52: joe_rgb=24'h524c43;
    8'h30: joe_rgb=24'h302921;
    8'h51: joe_rgb=24'h514c42;
    8'hd9: joe_rgb=24'hd9c4b3;
    8'hf6: joe_rgb=24'hf6e6d2;
    8'hd7: joe_rgb=24'hd7c2b1;
    8'h4e: joe_rgb=24'h4e4a40;
    8'h3c: joe_rgb=24'h3c352d;
    8'h34: joe_rgb=24'h34322c;
    8'heb: joe_rgb=24'hebe0d5;
    8'hea: joe_rgb=24'heae4d6;
    8'hca: joe_rgb=24'hcaa697;
    8'hd0: joe_rgb=24'hd0ac9d;
    8'hcf: joe_rgb=24'hcfaa9c;
    8'hd2: joe_rgb=24'hd2b1a8;
    8'hce: joe_rgb=24'hcea79f;
    8'h3a: joe_rgb=24'h3a3e48;
    8'h10: joe_rgb=24'h10111e;
    8'h39: joe_rgb=24'h393d47;
    8'he4: joe_rgb=24'he4d4d4;
    8'he1: joe_rgb=24'he1d2d1;
    8'h36: joe_rgb=24'h363b44;
    8'h1e: joe_rgb=24'h1e202c;
    8'h15: joe_rgb=24'h151d2b;
    8'h84: joe_rgb=24'h847374;
    8'hd8: joe_rgb=24'hd8c1b7;
    8'hcc: joe_rgb=24'hcca394;
    8'h2c: joe_rgb=24'h2c2f31;
    8'h01: joe_rgb=24'h010005;
    8'h2b: joe_rgb=24'h2b2e30;
    8'h28: joe_rgb=24'h282b2e;
    8'h04: joe_rgb=24'h040b12;
    8'h7b: joe_rgb=24'h7b6a63;
    8'he3: joe_rgb=24'he3d2c9;
    8'h98: joe_rgb=24'h988f8b;
    8'he7: joe_rgb=24'he7d6cd;
    8'he9: joe_rgb=24'he9d8cf;
    8'hdd: joe_rgb=24'hddc7be;
    8'hf4: joe_rgb=24'hf4efed;
    8'hc0: joe_rgb=24'hc09381;
    8'hdc: joe_rgb=24'hdca38c;
    8'h5f: joe_rgb=24'h5f6b42;
    8'h00: joe_rgb=24'h005d85;
    8'h16: joe_rgb=24'h16667e;
    8'h1c: joe_rgb=24'h1c6f89;
    8'h1b: joe_rgb=24'h1b6d86;
    8'h18: joe_rgb=24'h186982;
    8'h60: joe_rgb=24'h606b42;
    8'hcd: joe_rgb=24'hcda69d;
    8'h64: joe_rgb=24'h64785a;
    8'h0e: joe_rgb=24'h0e6d98;
    8'h29: joe_rgb=24'h297186;
    8'h26: joe_rgb=24'h267188;
    8'h65: joe_rgb=24'h65785a;
    8'h4a: joe_rgb=24'h4a756f;
    8'h42: joe_rgb=24'h427577;
    8'h23: joe_rgb=24'h23718d;
    8'h2a: joe_rgb=24'h2a7288;
    8'h43: joe_rgb=24'h437577;
    8'h4b: joe_rgb=24'h4b756f;
    8'h78: joe_rgb=24'h787c52;
    8'h13: joe_rgb=24'h136f97;
    8'h79: joe_rgb=24'h797d52;
    8'hbd: joe_rgb=24'hbd831c;
    8'h55: joe_rgb=24'h557768;
    8'h2e: joe_rgb=24'h2e7385;
    8'h1f: joe_rgb=24'h1f7091;
    8'h33: joe_rgb=24'h337381;
    8'h20: joe_rgb=24'h207090;
    8'hd3: joe_rgb=24'hd3b4a7;
    8'hbb: joe_rgb=24'hbb8a77;
    8'h32: joe_rgb=24'h327a89;
    8'h37: joe_rgb=24'h375e68;
    8'h25: joe_rgb=24'h255773;
    8'h24: joe_rgb=24'h245773;
    8'h50: joe_rgb=24'h504423;
    8'h5c: joe_rgb=24'h5c5335;
    8'h67: joe_rgb=24'h675d41;
    8'h69: joe_rgb=24'h696043;
    8'h68: joe_rgb=24'h685f42;
    8'h6b: joe_rgb=24'h6b6141;
    8'h2f: joe_rgb=24'h2f4054;
    8'h62: joe_rgb=24'h62583b;
    8'h0c: joe_rgb=24'h0c1b28;
    8'h19: joe_rgb=24'h192937;
    8'h1d: joe_rgb=24'h1d2c39;
    8'h2d: joe_rgb=24'h2d3d4b;
    8'h6e: joe_rgb=24'h6e767c;
    8'h09: joe_rgb=24'h09223e;
    8'h22: joe_rgb=24'h223b5a;
    8'h21: joe_rgb=24'h213a57;
    8'h05: joe_rgb=24'h051d39;
    8'h31: joe_rgb=24'h314556;
    8'h35: joe_rgb=24'h354555;
    8'h02: joe_rgb=24'h021728;
    8'h14: joe_rgb=24'h142b3b;
    8'h1a: joe_rgb=24'h1a2934;
    8'h77: joe_rgb=24'h777e82;
    8'h3b: joe_rgb=24'h3b414a;
    8'h3d: joe_rgb=24'h3d3030;
    8'h3f: joe_rgb=24'h3f3130;
    8'h47: joe_rgb=24'h47535d;
    8'h7c: joe_rgb=24'h7c8388;
    8'h5a: joe_rgb=24'h5a362a;
    8'h11: joe_rgb=24'h11212d;
    8'h40: joe_rgb=24'h40190c;
    8'h49: joe_rgb=24'h492215;
    8'h41: joe_rgb=24'h413f46;
    8'h3e: joe_rgb=24'h3e4e5e;
    8'h5d: joe_rgb=24'h5d666c;
    8'h57: joe_rgb=24'h573428;
    8'h56: joe_rgb=24'h563327;
    8'h58: joe_rgb=24'h583529;
    8'h12: joe_rgb=24'h122939;
    8'h4d: joe_rgb=24'h4d281c;
    8'h54: joe_rgb=24'h543227;
    8'h59: joe_rgb=24'h59372c;
    8'h63: joe_rgb=24'h63473c;
    8'h61: joe_rgb=24'h613e33;
    8'h53: joe_rgb=24'h533126;
    8'h27: joe_rgb=24'h273d4f;
    8'h4c: joe_rgb=24'h4c2418;
    8'h74: joe_rgb=24'h744f43;
    8'h48: joe_rgb=24'h483e3f;
    8'h38: joe_rgb=24'h384857;
    8'h70: joe_rgb=24'h704c40;
    8'h5e: joe_rgb=24'h5e382b;
    8'h03: joe_rgb=24'h031320;
    8'h73: joe_rgb=24'h734e42;
    8'h0f: joe_rgb=24'h0f1f2f;
    8'h72: joe_rgb=24'h724d41;
    8'h76: joe_rgb=24'h765145;
    8'h17: joe_rgb=24'h172736;
    8'h0a: joe_rgb=24'h0a1b2b;
    8'h75: joe_rgb=24'h755044;
    8'h0d: joe_rgb=24'h0d1e2d;
    8'h07: joe_rgb=24'h071929;
    8'h85: joe_rgb=24'h858c8f;
    8'h0b: joe_rgb=24'h0b1b2a;
    8'h4f: joe_rgb=24'h4f362f;
    8'h45: joe_rgb=24'h453a39;
    8'h44: joe_rgb=24'h441c0f;
    8'h86: joe_rgb=24'h868c8e;
    8'h6a: joe_rgb=24'h6a463b;
    8'h6c: joe_rgb=24'h6c483d;
    8'h6d: joe_rgb=24'h6d4c40;
    8'h7f: joe_rgb=24'h7f5b4f;

    default: joe_rgb=24'hffffff;
    endcase
    end
endmodule
