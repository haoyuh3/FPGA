`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/10/24 12:04:37
// Design Name: 
// Module Name: colormapper
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
// draw x and draw y is the current place use front to decide whether to draw
// x15  x,y-> 


module colormapper(input  logic [9:0] DrawX, DrawY,
                       output logic [3:0]  Red, Green, Blue

    );
    
endmodule
